
`timescale 1ns/1ns
module IM (input [31:0] address, output [31:0] instruction);

	parameter integer l = 500;
	reg [31:0] ins [1000:0];
	assign instruction = ins[address];

	initial begin
		for (int i = 0; i <= l; i++) begin
			ins[i] = 32'b0;
			// ins[i] = {6'b000001, 5'd1, 5'd1, 16'd255}; //addi R0, R1, 255
		end

		// ins[0] = {6'b000001, 5'd0, 5'd1, 16'd20}; // addi R0, R1, 40
		// ins[4] = {6'b000001, 5'd0, 5'd2, 16'd20}; // addi R0, R2, 20
		// ins[8] = {6'b000001, 5'd0, 5'd3, 16'd20}; // addi R0, R3, 40
		// ins[8] = {6'b000101, 5'd1, 5'd2, 16'd24}; // beq R1, R2, 16
		// ins[12] = {6'b000000, 5'd1, 5'd2, 5'd3, 6'b000001}; // sub R1, R2, R3

		// ins[16] = {6'b000101, 5'd2, 5'd3, 16'd32}; // beq R1, R2, 16

		// ins[8] = {6'b000100, 5'd2, 5'd1, 16'd0}; // sw R1, 0(R2)

		ins[0] = {6'b000000, 5'd0, 5'd0, 5'd4, 5'd0, 6'b000000}; // add R4, R0, R0
		ins[4] = {6'b000001, 5'd0, 5'd10, 16'd40}; // addi R0, R10, 40
		ins[8] = {6'b000101, 5'd4, 5'd10, 16'd32}; // beq R10, R4, 32
		ins[12] = {6'b000011, 5'd4, 5'd1, 16'd1000}; // lw R1, 1000(R4)
		ins[16] = {6'b000011, 5'd4, 5'd2, 16'd2000}; // lw R2, 2000(R4)
		ins[20] = {6'b000000, 5'd1, 5'd2, 5'd3, 5'd0, 6'b000000}; // add R3, R1, R2
		ins[24] = {6'b000100, 5'd4, 5'd3, 16'd3000}; // sw R3, 3000(R4)
		ins[28] = {6'b000001, 5'd4, 5'd4, 16'd4}; // addi R4, R4, 4
		ins[32] = {6'b000111, 26'd2}; // j 8 // j 2<<2

		ins[100] = {6'b000001, 5'd0, 5'd1, 16'd1}; // addi R1, R0, 1

		ins[104] = {6'b000001, 5'd0, 5'd4, 16'd1000}; // addi R4, R0, 1000
		ins[108] = {6'b000000, 5'd0, 5'd0, 5'd5, 5'd0, 6'b000000};// add R5, R0, R0

		ins[112] = {6'b000001, 5'd0, 5'd6, 16'd80};// addi R6, R0, 80

		ins[116] = {6'b000011, 5'd0, 5'd10, 16'd1000};// lw R10, 1000(R0)
		ins[120] = {6'b000000, 5'd0, 5'd0, 5'd11, 5'd0, 6'b000000}; // add R11, R0, R0
		ins[124] = {6'b000101, 5'd5, 5'd6, 16'd32}; // beq R5, R6, 32
		ins[128] = {6'b000011, 5'd5, 5'd12, 16'd1000};// lw R12, 1000(R5)
		ins[132] = {6'b000000, 5'd12, 5'd10, 5'd13, 5'd0, 6'b001000};// slt R13, R12, R10
		ins[136] = {6'b000101, 5'd1, 5'd13, 16'd8};  // beq R1, R13, 8
	
		ins[140] = {6'b000001, 5'd4, 5'd4, 16'd4};// addi R4, R4, 4
		ins[144] = {6'b000001, 5'd5, 5'd5, 16'd4};// addi R5, R5, 4
		ins[148] = {6'b000000, 5'd0, 5'd12, 5'd10, 5'd0, 6'b000000};// add R10, R12, R0
		ins[152] = {6'b000000, 5'd0, 5'd4, 5'd11, 5'd0, 6'b000000};// add R11, R4, R0

		ins[156] = {6'b000111, 26'd31}; // j 124 // j 6<<2

		ins[160] = {6'b000100, 5'd0, 5'd10, 16'd2000}; // sw R10, 2000(R0)
		ins[164] = {6'b000100, 5'd0, 5'd11, 16'd2004};// sw R11, 2004(R0) 

	end;
endmodule	


