
// module ErrorDP(input clk, rst, input [19:0] x, y, B0, B1, output [19:0] E);
//     wire [19:0] B1x, ysubB0;
//     Multiplier mulb1x(x, B1, B1x);
//     AddOrSub subyb0(y, B0, 0, ysubB0);
//     AddOrSub subyb0(ysubB0, B1x, 0, E);
//     Register20bit regE(clk, rst)
// endmodule
