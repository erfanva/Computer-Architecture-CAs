
module DataLoaderDP(input clk, rst);

endmodule