
module DataLoaderCU(input clk, rst);
    
endmodule